module memory (clk, addr);
	input clk;
	input[28:0] addr;
	reg[31:0] Mem[(1<<28)-1];
	always @(posedge clk) begin
		
	/*
		Mem[0] = 28'b 0000000000000000000000000000;
		Mem[1] = 28'b 0000000000000000000000000001;
		Mem[2] = 28'b 0000000000000000000000000010;
		Mem[3] = 28'b 0000000000000000000000000011;
		Mem[4] = 28'b 0000000000000000000000000100;
		Mem[5] = 28'b 0000000000000000000000000101;
		Mem[6] = 28'b 0000000000000000000000000110;
		Mem[7] = 28'b 0000000000000000000000000111;
		Mem[8] = 28'b 0000000000000000000000001000;
		Mem[9] = 28'b 0000000000000000000000001001;
		Mem[10] = 28'b 0000000000000000000000001010;
		Mem[11] = 28'b 0000000000000000000000001011;
		Mem[12] = 28'b 0000000000000000000000001100;
		Mem[13] = 28'b 0000000000000000000000001101;
		Mem[14] = 28'b 0000000000000000000000001110;
		Mem[15] = 28'b 0000000000000000000000001111;
		Mem[16] = 28'b 0000000000000000000000000000;
		Mem[17] = 28'b 0000000000000000000000000001;
		Mem[18] = 28'b 0000000000000000000000000010;
		Mem[19] = 28'b 0000000000000000000000000011;
		Mem[20] = 28'b 0000000000000000000000000100;
		Mem[21] = 28'b 0000000000000000000000000101;
		Mem[22] = 28'b 0000000000000000000000000110;
		Mem[23] = 28'b 0000000000000000000000000111;
		Mem[24] = 28'b 0000000000000000000000001000;
		Mem[25] = 28'b 0000000000000000000000001001;
		Mem[26] = 28'b 0000000000000000000000001010;
		Mem[27] = 28'b 0000000000000000000000001011;
		Mem[28] = 28'b 0000000000000000000000001100;
		Mem[29] = 28'b 0000000000000000000000001101;
		Mem[30] = 28'b 0000000000000000000000001110;
		Mem[31] = 28'b 0000000000000000000000001111;
		Mem[32] = 28'b 0000000000000000000000000000;
		Mem[33] = 28'b 0000000000000000000000000001;
		Mem[34] = 28'b 0000000000000000000000000010;
		Mem[35] = 28'b 0000000000000000000000000011;
		Mem[36] = 28'b 0000000000000000000000000100;
		Mem[37] = 28'b 0000000000000000000000000101;
		Mem[38] = 28'b 0000000000000000000000000110;
		Mem[39] = 28'b 0000000000000000000000000111;
		Mem[40] = 28'b 0000000000000000000000001000;
		Mem[41] = 28'b 0000000000000000000000001001;
		Mem[42] = 28'b 0000000000000000000000001010;
		Mem[43] = 28'b 0000000000000000000000001011;
		Mem[44] = 28'b 0000000000000000000000001100;
		Mem[45] = 28'b 0000000000000000000000001101;
		Mem[46] = 28'b 0000000000000000000000001110;
		Mem[47] = 28'b 0000000000000000000000001111;
		Mem[48] = 28'b 0000000000000000000000000000;
		Mem[49] = 28'b 0000000000000000000000000001;
		Mem[50] = 28'b 0000000000000000000000000010;
		Mem[51] = 28'b 0000000000000000000000000011;
		Mem[52] = 28'b 0000000000000000000000000100;
		Mem[53] = 28'b 0000000000000000000000000101;
		Mem[54] = 28'b 0000000000000000000000000110;
		Mem[55] = 28'b 0000000000000000000000000111;
		Mem[56] = 28'b 0000000000000000000000001000;
		Mem[57] = 28'b 0000000000000000000000001001;
		Mem[58] = 28'b 0000000000000000000000001010;
		Mem[59] = 28'b 0000000000000000000000001011;
		Mem[60] = 28'b 0000000000000000000000001100;
		Mem[61] = 28'b 0000000000000000000000001101;
		Mem[62] = 28'b 0000000000000000000000001110;
		Mem[63] = 28'b 0000000000000000000000001111;

		Mem[64] = 28'b 0000000000000000000000000000;
		Mem[65] = 28'b 0000000000000000000000000001;
		Mem[66] = 28'b 0000000000000000000000000010;
		Mem[67] = 28'b 0000000000000000000000000011;
		Mem[68] = 28'b 0000000000000000000000000100;
		Mem[69] = 28'b 0000000000000000000000000101;
		Mem[70] = 28'b 0000000000000000000000000110;
		Mem[71] = 28'b 0000000000000000000000000111;
		Mem[72] = 28'b 0000000000000000000000001000;
		Mem[73] = 28'b 0000000000000000000000001001;
		Mem[74] = 28'b 0000000000000000000000001010;
		Mem[75] = 28'b 0000000000000000000000001011;
		Mem[76] = 28'b 0000000000000000000000001100;
		Mem[77] = 28'b 0000000000000000000000001101;
		Mem[78] = 28'b 0000000000000000000000001110;
		Mem[79] = 28'b 0000000000000000000000001111;
		Mem[80] = 28'b 0000000000000000000000000000;
		Mem[81] = 28'b 0000000000000000000000000001;
		Mem[82] = 28'b 0000000000000000000000000010;
		Mem[83] = 28'b 0000000000000000000000000011;
		Mem[84] = 28'b 0000000000000000000000000100;
		Mem[85] = 28'b 0000000000000000000000000101;
		Mem[86] = 28'b 0000000000000000000000000110;
		Mem[87] = 28'b 0000000000000000000000000111;
		Mem[88] = 28'b 0000000000000000000000001000;
		Mem[89] = 28'b 0000000000000000000000001001;
		Mem[90] = 28'b 0000000000000000000000001010;
		Mem[91] = 28'b 0000000000000000000000001011;
		Mem[92] = 28'b 0000000000000000000000001100;
		Mem[93] = 28'b 0000000000000000000000001101;
		Mem[94] = 28'b 0000000000000000000000001110;
		Mem[95] = 28'b 0000000000000000000000001111;
		Mem[96] = 28'b 0000000000000000000000000000;
		Mem[97] = 28'b 0000000000000000000000000001;
		Mem[98] = 28'b 0000000000000000000000000010;
		Mem[99] = 28'b 0000000000000000000000000011;
		Mem[100] = 28'b 0000000000000000000000000100;
		Mem[101] = 28'b 0000000000000000000000000101;
		Mem[102] = 28'b 0000000000000000000000000110;
		Mem[103] = 28'b 0000000000000000000000000111;
		Mem[104] = 28'b 0000000000000000000000001000;
		Mem[105] = 28'b 0000000000000000000000001001;
		Mem[106] = 28'b 0000000000000000000000001010;
		Mem[107] = 28'b 0000000000000000000000001011;
		Mem[108] = 28'b 0000000000000000000000001100;
		Mem[109] = 28'b 0000000000000000000000001101;
		Mem[110] = 28'b 0000000000000000000000001110;
		Mem[111] = 28'b 0000000000000000000000001111;
		Mem[112] = 28'b 0000000000000000000000000000;
		Mem[113] = 28'b 0000000000000000000000000001;
		Mem[114] = 28'b 0000000000000000000000000010;
		Mem[115] = 28'b 0000000000000000000000000011;
		Mem[116] = 28'b 0000000000000000000000000100;
		Mem[117] = 28'b 0000000000000000000000000101;
		Mem[118] = 28'b 0000000000000000000000000110;
		Mem[119] = 28'b 0000000000000000000000000111;
		Mem[120] = 28'b 0000000000000000000000001000;
		Mem[121] = 28'b 0000000000000000000000001001;
		Mem[122] = 28'b 0000000000000000000000001010;
		Mem[123] = 28'b 0000000000000000000000001011;
		Mem[124] = 28'b 0000000000000000000000001100;
		Mem[125] = 28'b 0000000000000000000000001101;
		Mem[126] = 28'b 0000000000000000000000001110;
		Mem[127] = 28'b 0000000000000000000000001111;
		*/
	end
endmodule


